module chip (
    inout  [2:0] P_GPIO,
    // RF I/O Pins
    input  P_RF_RX,
    output P_RF_TX,
    inout  [4:1] P_ANALOG_TEST,
    // CPU I/O Pins,
    output P_UART_TX,
    input  P_UART_RX,
    input  P_MSEL,
    input  P_JTAG_TCK,
    output P_JTAG_TDO,
    input  P_JTAG_TMS,
    input  P_JTAG_TDI,
    output P_SPI_CS,
    output P_SPI_SCK,
    input  [3:0] P_SPI_DQ,
    output P_TL_CLK,
    input  P_TL_IN_DAT,
    output P_TL_IN_RDY,
    input  P_TL_IN_VAL,
    output P_TL_OUT_DAT,
    input  P_TL_OUT_RDY,
    output P_TL_OUT_VAL,
    //DBB I/O Pin,
    output P_DBB_OFF_CHIP_MODE_TX,
    output P_DBB_OFF_CHIP_MODE_RX,
    // Power/Clocking I/O Pins,
    input  P_RESET,
    input  P_CPU_REF_CLK,
    input  P_RF_REF_CLK,
    input  P_V_BAT,
    input  P_V_REF,
    input  P_I_REF,
    input  P_GND,
    input  P_IO_PWR,
    input  P_LDO_EN,
    input  P_VDD_D,
    input  P_VDD_A
);
    
    //GPIO and Analog
    wire [2:0] gpio_rd_d, gpio_wr_d, gpio_wr_enn;
    wire [3:0] spi_dq_rd_d, spi_dq_wr_d, spi_dq_wr_enn;
    //Digital
    wire uart_tx, uart_rx, msel, jtag_tck, jtag_tdo_data, jtag_tdo_driven, jtag_tms, jtag_tdi, spi_cs, spi_sck ,spi_dq_0, spi_dq_1, spi_dq_2, spi_dq_3, tl_clk, tl_in_dat, tl_in_rdy, tl_in_val, tl_out_dat, tl_out_rdy, tl_out_val;
    //DBB and Power
    wire dbb_off_chip_mode_tx, dbb_off_chip_mode_rx, reset, cpu_ref_clk, clk_over;

    core core(
        .gpio_rd_d(gpio_rd_d),
        .gpio_wr_d(gpio_wr_d),
        .gpio_wr_enn(gpio_wr_enn),
    // RF I/O Pins
        .rf_rx(P_RF_RX),
        .rf_tx(P_RF_TX),
        .analog_test(P_ANALOG_TEST),
    // CPU I/O Pins,
        .uart_tx(uart_tx),
        .uart_rx(uart_rx),
        .msel(msel),
        .jtag_tck(jtag_tck),
        .jtag_tdo_data(jtag_tdo_data),
        .jtag_tdo_driven(jtag_tdo_driven),
        .jtag_tms(jtag_tms),
        .jtag_tdi(jtag_tdi),
        .spi_cs(spi_cs),
        .spi_sck(spi_sck),
        .spi_dq_rd_d(spi_dq_rd_d),
        .spi_dq_wr_d(spi_dq_wr_d),
        .spi_dq_wr_enn(spi_dq_wr_enn),
        .tl_clk(tl_clk),
        .tl_in_dat(tl_in_dat),
        .tl_in_rdy(tl_in_rdy),
        .tl_in_val(tl_in_val),
        .tl_out_dat(tl_out_dat),
        .tl_out_rdy(tl_out_rdy),
        .tl_out_val(tl_out_val),
    //DBB I/O Pin,
        .dbb_off_chip_mode_tx(dbb_off_chip_mode_tx),
        .dbb_off_chip_mode_rx(dbb_off_chip_mode_rx),
    // Power/Clocking I/O Pins,
        .reset(reset),
        .cpu_ref_clk(cpu_ref_clk),
        .rf_ref_clk(P_RF_REF_CLK),
        .v_bat(P_V_BAT),
        .v_ref(P_V_REF),
        .i_ref(P_I_REF),
        .gnd(P_GND),
        .io_pwr(P_IO_PWR),
        .ldo_en(P_LDO_EN),
        .vdd_d(P_VDD_D),
        .vdd_a(P_VDD_A)
    );
    
    io_ring_clamped IoRing(
        .gpio_rd_d(gpio_rd_d),
        .gpio_wr_d(gpio_wr_d),
        .gpio_wr_enn(gpio_wr_enn),
    // CPU I/O Pins,
        .uart_tx(uart_tx),
        .uart_rx(uart_rx),
        .msel(msel),
        .jtag_tck(jtag_tck),
        .jtag_tdo(jtag_tdo_data),
        .jtag_tdo_driven(jtag_tdo_driven),
        .jtag_tms(jtag_tms),
        .jtag_tdi(jtag_tdi),
        .spi_cs(spi_cs),
        .spi_sck(spi_sck),
        .spi_dq_rd_d(spi_dq_rd_d),
        .spi_dq_wr_d(spi_dq_wr_d),
        .spi_dq_wr_enn(spi_dq_wr_enn),
        .tl_clk(tl_clk),
        .tl_in_dat(tl_in_dat),
        .tl_in_rdy(tl_in_rdy),
        .tl_in_val(tl_in_val),
        .tl_out_dat(tl_out_dat),
        .tl_out_rdy(tl_out_rdy),
        .tl_out_val(tl_out_val),
    //DBB I/O Pin,
        .dbb_off_chip_mode_tx(dbb_off_chip_mode_tx),
        .dbb_off_chip_mode_rx(dbb_off_chip_mode_rx),
    // Power/Clocking I/O Pins,
        .reset(reset),
        .cpu_ref_clk(cpu_ref_clk),
    /*************IO_Ring to Pad_Ring***************/
        .P_GPIO(P_GPIO),
    // RF I/O Pins
        .P_RF_RX(P_RF_RX),
        .P_RF_TX(P_RF_TX),
        .P_ANALOG_TEST_1(P_ANALOG_TEST[1]),
        .P_ANALOG_TEST_2(P_ANALOG_TEST[2]),
        .P_ANALOG_TEST_3(P_ANALOG_TEST[3]),
        .P_ANALOG_TEST_4(P_ANALOG_TEST[4]),
    // CPU I/O Pins,
        .P_UART_TX(P_UART_TX),
        .P_UART_RX(P_UART_RX),
        .P_MSEL(P_MSEL),
        .P_JTAG_TCK(P_JTAG_TCK),
        .P_JTAG_TDO(P_JTAG_TDO),
        .P_JTAG_TMS(P_JTAG_TMS),
        .P_JTAG_TDI(P_JTAG_TDI),
        .P_SPI_CS(P_SPI_CS),
        .P_SPI_SCK(P_SPI_SCK),
        .P_SPI_DQ(P_SPI_DQ),
        .P_TL_CLK(P_TL_CLK),
        .P_TL_IN_DAT(P_TL_IN_DAT),
        .P_TL_IN_RDY(P_TL_IN_RDY),
        .P_TL_IN_VAL(P_TL_IN_VAL),
        .P_TL_OUT_DAT(P_TL_OUT_DAT),
        .P_TL_OUT_RDY(P_TL_OUT_RDY),
        .P_TL_OUT_VAL(P_TL_OUT_VAL),
    //DBB I/O Pin,
        .P_DBB_OFF_CHIP_MODE_TX(P_DBB_OFF_CHIP_MODE_TX),
        .P_DBB_OFF_CHIP_MODE_RX(P_DBB_OFF_CHIP_MODE_RX),
    // Power/Clocking I/O Pins,
        .P_RESET(P_RESET),
        .P_CPU_REF_CLK(P_CPU_REF_CLK),
        .P_RF_REF_CLK(P_RF_REF_CLK),
        .P_V_BAT(P_V_BAT),
        .P_V_REF(P_V_REF),
        .P_I_REF(P_I_REF),
        .P_GND(P_GND),
        .P_IO_PWR(P_IO_PWR),
        .P_LDO_EN(P_LDO_EN),
        .P_VDD_D(P_VDD_D),
        .P_VDD_A(P_VDD_A)
    );

endmodule
