module ChipTop( // @[chipyard.TestHarness.EE290CBLEConfig.fir 261941:2]
  input         jtag_TCK, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295019:4]
  input         jtag_TMS, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295019:4]
  input         jtag_TDI, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295019:4]
  output        jtag_TDO_data, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295019:4]
  output        jtag_TDO_driven, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295019:4]
  output        serial_tl_clock, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  output        serial_tl_bits_in_ready, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  input         serial_tl_bits_in_valid, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  input         serial_tl_bits_in_bits, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  input         serial_tl_bits_out_ready, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  output        serial_tl_bits_out_valid, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  output        serial_tl_bits_out_bits, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295020:4]
  output        baseband_offChipMode_rx, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output        baseband_offChipMode_tx, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_data_tx_loFSK, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  input  [7:0]  baseband_data_rx_i_data, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  input  [7:0]  baseband_data_rx_q_data, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_data_loCT, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [10:0] baseband_data_pllD, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g4, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g5, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g6, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [7:0]  baseband_tuning_trim_g7, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_mixer_r0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_mixer_r1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_mixer_r2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_mixer_r3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [9:0]  baseband_tuning_i_vgaAtten, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r4, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r5, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r6, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r7, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r8, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_i_filter_r9, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [9:0]  baseband_tuning_q_vgaAtten, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r4, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r5, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r6, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r7, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r8, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [3:0]  baseband_tuning_q_filter_r9, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [5:0]  baseband_tuning_dac_t0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [5:0]  baseband_tuning_dac_t1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [5:0]  baseband_tuning_dac_t2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [5:0]  baseband_tuning_dac_t3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [4:0]  baseband_tuning_enable_rx_i, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [4:0]  baseband_tuning_enable_rx_q, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output        baseband_tuning_enable_debug, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [9:0]  baseband_tuning_mux_dbg_in, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  output [9:0]  baseband_tuning_mux_dbg_out, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295021:4]
  inout         gpio_0_0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295022:4]
  inout         gpio_0_1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295023:4]
  output        spi_0_sck, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  output        spi_0_cs_0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  inout         spi_0_dq_0, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  inout         spi_0_dq_1, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  inout         spi_0_dq_2, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  inout         spi_0_dq_3, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295024:4]
  output        uart_0_txd, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295025:4]
  input         uart_0_rxd, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295025:4]
  input         bsel, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295026:4]
  input         reset_wire_reset, // @[chipyard.TestHarness.EE290CBLEConfig.fir 295027:4]
  input         clock // @[chipyard.TestHarness.EE290CBLEConfig.fir 295028:4]
);
endmodule 
