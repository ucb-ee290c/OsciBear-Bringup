module rf_top(
       inout VDDA,
       inout VSS,
       inout rf_ref_clk,
       inout cpu_clk,
       inout pll_cref,
       inout lo_cref,
       inout div_cref,
       inout bp_cref_i,
       inout bp_cref_q,
       inout vga_cref_0i,
       inout vga_cref_1i,
       inout vga_cref_0q,
       inout vga_cref_1q,
       inout mixer_cref,
       inout buff_cref_i,
       inout buff_cref_q,
       inout test_cref,
       inout analog_test1,
       inout analog_test2,
       inout analog_test3,
       inout analog_test4,
       inout test_en,
       inout rf_clk_sel,
       inout analog_test2_sel,
       inout [9:0] mux_dbg_in,
       inout [9:0] mux_dbg_out,
       inout [7:0] i_adc_code,     
       inout [7:0] q_adc_code, 
       inout i_adc_data_valid,
       inout q_adc_data_valid,
       inout [4:0] i_enable,
       inout [4:0] q_enable,
       inout RF_TX,
       inout RF_IN,
       inout [7:0] lo_fsk_tune,
       inout [5:0] lo_coarse_tune,
       inout [10:0] pll_div,
       inout cc_enable, 
       inout ref_sel, 
       inout pll_sign, 
       inout [5:0] pll_idac,
       inout lo_enable,
       inout [3:0] filter_res0i,
       inout [3:0] filter_res1i, 
       inout [3:0] filter_res2i,
       inout [3:0] filter_res3i,
       inout [3:0] filter_res4i,
       inout [3:0] filter_res5i,
       inout [3:0] filter_res6i,
       inout [3:0] filter_res7i,
       inout [3:0] filter_res8i,
       inout [3:0] filter_res9i,
       inout [3:0] filter_res0q,
       inout [3:0] filter_res1q, 
       inout [3:0] filter_res2q,
       inout [3:0] filter_res3q,
       inout [3:0] filter_res4q,
       inout [3:0] filter_res5q,
       inout [3:0] filter_res6q,
       inout [3:0] filter_res7q,
       inout [3:0] filter_res8q,
       inout [3:0] filter_res9q,
       inout [9:0] VGA_atteni, 
       inout [9:0] VGA_attenq, 
       inout [5:0] current_dac_0i,
       inout [5:0] current_dac_1i,
       inout [5:0] current_dac_0q,
       inout [5:0] current_dac_1q,
       inout [3:0] mix_res_in,
       inout [3:0] mix_res_ip,
       inout [3:0] mix_res_qn,
       inout [3:0] mix_res_qp
    );

endmodule
