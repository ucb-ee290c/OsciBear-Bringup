//This will be the pad ring
module io_ring (
/*************chip_top io_ring***************/
    inout gpio_0,
    inout gpio_1,
    inout gpio_2,
// RF I/O Pins
    input rf_rx,
    output rf_tx,
    inout analog_test_1,
    inout analog_test_2,
    inout analog_test_3,
    inout analog_test_4, 
// CPU I/O Pins,
    output uart_tx,
    input uart_rx,
    input msel,
    input jtag_tck,
    output jtag_tdo,
    input jtag_tms,
    input jtag_tdi,
    output spi_cs,
    output spi_sck,
    input spi_dq_0,
    input spi_dq_1,
    input spi_dq_2,
    input spi_dq_3,
    output tl_clk,
    input tl_in_dat,
    output tl_in_rdy,
    input tl_in_val,
    output tl_out_dat,
    input tl_out_rdy,
    output tl_out_val,
//DBB I/O Pin,
    output dbb_off_chip_mode_tx,
    output dbb_off_chip_mode_rx,
// Power/Clocking I/O Pins,
    input reset,
    input cpu_ref_clk,
    input rf_ref_clk,
    input v_bat,
    input v_ref,
    input i_ref,
    input gnd,
    input io_pwr,
    input ldo_en,
    input vdd_d,
    input vdd_a,

/*************IO_Ring to Pad_Ring***************/
    inout GPIO_0,
    inout GPIO_1,
    inout GPIO_2,
// RF I/O Pins
    input RF_RX,
    output RF_TX,
    inout ANALOG_TEST_1,
    inout ANALOG_TEST_2,
    inout ANALOG_TEST_3,
    inout ANALOG_TEST_4, 
// CPU I/O Pins,
    output UART_TX,
    input UART_RX,
    input MSEL,
    input JTAG_TCK,
    output JTAG_TDO,
    input JTAG_TMS,
    input JTAG_TDI,
    output SPI_CS,
    output SPI_SCK,
    input SPI_DQ_0,
    input SPI_DQ_1,
    input SPI_DQ_2,
    input SPI_DQ_3,
    output TL_CLK,
    input TL_IN_DAT,
    output TL_IN_RDY,
    input TL_IN_VAL,
    output TL_OUT_DAT,
    input TL_OUT_RDY,
    output TL_OUT_VAL,
//DBB I/O Pin,
    output DBB_OFF_CHIP_MODE_TX,
    output DBB_OFF_CHIP_MODE_RX,
// Power/Clocking I/O Pins,
    input RESET,
    input CPU_REF_CLK,
    input RF_REF_CLK,
    input V_BAT,
    input V_REF,
    input I_REF,
    input GND_0,
    input GND_1,
    input GND_2,
    input GND_3,
    input GND_4,
    input GND_5,
    input GND_6,
    input IO_PWR,
    input LDO_EN,
    input VDD_D,
    input VDD_A
);

